`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    15:51:41 08/31/2011 
// Design Name: 
// Module Name:    ALUmod 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module ALUmod(
    input [15:0] A,
    input [15:0] B,
    input [3:0] opcode,
    output [15:0] S,
    input [3:0] opext,
    output [4:0] CLFZN
    );

//start always block and add all the different executions

always@(A,B,opcode)
	begin
	
	
	
	end


endmodule
