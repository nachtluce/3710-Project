`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    16:40:37 10/06/2011 
// Design Name: 
// Module Name:    bitGen_minimum 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module bitGen_minimum(
    input bright,
    input [9:0] hCount,
    input [9:0] vCount,
    output [2:0] rgb
    );


endmodule
